
 ////////////////////////////////////////////////////////////////////////
 //devloper name : 
 //date   : 
 //Description : 
 //////////////////////////////////////////////////////////////////////

 class axi_slave_env_config extends uvm_object;

 ////////////////////////////////////////////////////////////////////////
 //Method name : 
 //Arguments   :  
 //Description : 
 //////////////////////////////////////////////////////////////////////
 
 function new(string str = "axi_slave_env_config"); 
    super.new(str);
 endfunction : new


//for enabling coverage checker and scoreboard pins
 bit coverage_pin;
 bit scoreboard_pin;
 bit checker_pin;

 endclass
 









