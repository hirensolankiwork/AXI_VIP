
////////////////////////////////////////////////////////////////////////
//devloper name : siddharth 
//date   :  24/07/2023
//Description : 
//////////////////////////////////////////////////////////////////////

class slave_sequencer extends uvm_sequencer#(axi_slave_seq_item);
 `uvm_component_utils(slave_sequencer)
  bit[7:0] slv_mem[int];
  int len[];
  axi_slave_seq_item  tr_h;
  virtual axi_interface axi_inf;
  uvm_blocking_get_port #(axi_slave_seq_item) get_port;
  
  ////////////////////////////////////////////////////////////////////////
  //Method name : 
  //Arguments   :  
  //Description : 
  //////////////////////////////////////////////////////////////////////
  function new(string str = "slave_sequencer",uvm_component parent = null);
    super.new(str,parent);
    tr_h = new();
    get_port = new("get_port",this);
  endfunction
  ////////////////////////////////////////////////////////////////////////
  //Method name : 
  //Arguments   :  
  //Description : 
  /////////////////////////////////////////////////////////////////////
endclass
